LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BTN_COUNTER IS
  PORT(
  CLK_IN:IN STD_LOGIC;
  EN_IN:IN STD_LOGIC;
  STATE_OUT:BUFFER STD_LOGIC
  );
END ENTITY BTN_COUNTER;

ARCHITECTURE BEHAVE OF BTN_COUNTER IS
SIGNAL COUNT:INTEGER RANGE 0 TO 3;
BEGIN
  PROCESS(CLK_IN)
  BEGIN
    IF CLK_IN'EVENT AND CLK_IN='0' THEN
	    IF EN_IN='1' THEN
		    IF COUNT>= 3  THEN
			    STATE_OUT<='1';
			 ELSE
			    COUNT<=COUNT+1;
			 END IF;
		 ELSE
		    STATE_OUT<='0';
			 COUNT<=0;
		 END IF;
	 END IF;
  END PROCESS;
END BEHAVE;