LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--行信号读值，列信号循环写0
ENTITY BTN_DETECT IS
  PORT(
  CLK_IN:IN STD_LOGIC;
--  ROW0_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
--  ROW1_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
--  ROW2_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
--  ROW3_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
  KBROW:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0);
  KBCOL0:IN STD_LOGIC;
  KBCOL1:IN STD_LOGIC;
  KBCOL2:IN STD_LOGIC;
  KBCOL3:IN STD_LOGIC
  );
END ENTITY BTN_DETECT;

ARCHITECTURE DETECTION OF BTN_DETECT IS
SIGNAL COUNT:INTEGER RANGE 0 TO 3;
BEGIN
  CLK_COUNT:PROCESS(CLK_IN)
  BEGIN
    IF CLK_IN'EVENT AND CLK_IN='0' THEN
	   IF COUNT=3 THEN
		   COUNT<=0;
		ELSE
	      COUNT<=COUNT+1;
		END IF;	
	 END IF;
  END PROCESS CLK_COUNT;
  
  SCAN:PROCESS(COUNT,KBCOL0,KBCOL1,KBCOL2,KBCOL3)
  BEGIN
    CASE COUNT IS
	   WHEN 0 =>
		  IF KBCOL0='1' THEN KBROW(0)<='1'; ELSE KBROW(0)<='0'; END IF;
		  IF KBCOL1='1' THEN KBROW(1)<='1'; ELSE KBROW(1)<='0'; END IF;
		  IF KBCOL2='1' THEN KBROW(2)<='1'; ELSE KBROW(2)<='0'; END IF;
		  IF KBCOL3='1' THEN KBROW(3)<='1'; ELSE KBROW(3)<='0'; END IF;
		WHEN 1 =>
		  IF KBCOL0='1' THEN KBROW(0)<='1'; ELSE KBROW(0)<='0'; END IF;
		  IF KBCOL1='1' THEN KBROW(1)<='1'; ELSE KBROW(1)<='0'; END IF;
		  IF KBCOL2='1' THEN KBROW(2)<='1'; ELSE KBROW(2)<='0'; END IF;
		  IF KBCOL3='1' THEN KBROW(3)<='1'; ELSE KBROW(3)<='0'; END IF;
		WHEN 2 =>
		  IF KBCOL0='1' THEN KBROW(0)<='1'; ELSE KBROW(0)<='0'; END IF;
		  IF KBCOL1='1' THEN KBROW(1)<='1'; ELSE KBROW(1)<='0'; END IF;
		  IF KBCOL2='1' THEN KBROW(2)<='1'; ELSE KBROW(2)<='0'; END IF;
		  IF KBCOL3='1' THEN KBROW(3)<='1'; ELSE KBROW(3)<='0'; END IF;
		WHEN 3 =>
		  IF KBCOL0='1' THEN KBROW(0)<='1'; ELSE KBROW(0)<='0'; END IF;
		  IF KBCOL1='1' THEN KBROW(1)<='1'; ELSE KBROW(1)<='0'; END IF;
		  IF KBCOL2='1' THEN KBROW(2)<='1'; ELSE KBROW(2)<='0'; END IF;
		  IF KBCOL3='1' THEN KBROW(3)<='1'; ELSE KBROW(3)<='0'; END IF;	  
--	   WHEN 0 =>
--		  IF KBCOL0='1' THEN ROW0_OUT(0)<='1'; ELSE ROW0_OUT(0)<='0'; END IF;
--		  IF KBCOL1='1' THEN ROW0_OUT(1)<='1'; ELSE ROW0_OUT(1)<='0'; END IF;
--		  IF KBCOL2='1' THEN ROW0_OUT(2)<='1'; ELSE ROW0_OUT(2)<='0'; END IF;
--		  IF KBCOL3='1' THEN ROW0_OUT(3)<='1'; ELSE ROW0_OUT(3)<='0'; END IF;
--		WHEN 1 =>
--		  IF KBCOL0='1' THEN ROW1_OUT(0)<='1'; ELSE ROW1_OUT(0)<='0'; END IF;
--		  IF KBCOL1='1' THEN ROW1_OUT(1)<='1'; ELSE ROW1_OUT(1)<='0'; END IF;
--		  IF KBCOL2='1' THEN ROW1_OUT(2)<='1'; ELSE ROW1_OUT(2)<='0'; END IF;
--		  IF KBCOL3='1' THEN ROW1_OUT(3)<='1'; ELSE ROW1_OUT(3)<='0'; END IF;
--		WHEN 2 =>
--		  IF KBCOL0='1' THEN ROW2_OUT(0)<='1'; ELSE ROW2_OUT(0)<='0'; END IF;
--		  IF KBCOL1='1' THEN ROW2_OUT(1)<='1'; ELSE ROW2_OUT(1)<='0'; END IF;
--		  IF KBCOL2='1' THEN ROW2_OUT(2)<='1'; ELSE ROW2_OUT(2)<='0'; END IF;
--		  IF KBCOL3='1' THEN ROW2_OUT(3)<='1'; ELSE ROW2_OUT(3)<='0'; END IF;
--		WHEN 3 =>
--		  IF KBCOL0='1' THEN ROW3_OUT(0)<='1'; ELSE ROW3_OUT(0)<='0'; END IF;
--		  IF KBCOL1='1' THEN ROW3_OUT(1)<='1'; ELSE ROW3_OUT(1)<='0'; END IF;
--		  IF KBCOL2='1' THEN ROW3_OUT(2)<='1'; ELSE ROW3_OUT(2)<='0'; END IF;
--		  IF KBCOL3='1' THEN ROW3_OUT(3)<='1'; ELSE ROW3_OUT(3)<='0'; END IF;
	 END CASE;
  END PROCESS SCAN;
  
END DETECTION;
