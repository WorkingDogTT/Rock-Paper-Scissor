LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY DIVIDER_SERIAL IS
  PORT(
  CLK_IN    : IN STD_LOGIC;         --1kHz input clock
  CLK_512Hz : BUFFER STD_LOGIC;     --2x diff
  CLK_64Hz  : BUFFER STD_LOGIC;     --16x diff
  CLK_8Hz   : BUFFER STD_LOGIC;     --128x diff
  CLK_1Hz   : BUFFER STD_LOGIC      --1024x diff
  );
END DIVIDER_SERIAL;


ARCHITECTURE DIVIDE_SERIAL OF DIVIDER_SERIAL IS
--SIGNAL COUNT:INTEGER;
--SIGNAL COUNT_MAX:INTEGER;
  SIGNAL COUNT_1 : INTEGER RANGE 0 TO 3;
  SIGNAL COUNT_2 : INTEGER RANGE 0 TO 3;
  SIGNAL COUNT_3 : INTEGER RANGE 0 TO 3;
  
BEGIN

  PROCESS(CLK_IN)
  BEGIN
    IF (CLK_IN'EVENT AND CLK_IN='0') THEN
			 CLK_512Hz <= NOT CLK_512Hz;
	 END IF;
  END PROCESS; 
  
  PROCESS(CLK_512Hz)
  BEGIN
    IF (CLK_512Hz'EVENT AND CLK_512Hz='0') THEN
			 COUNT_1 <= COUNT_1+1;
			 IF (COUNT_1 = 3) THEN
			   COUNT_1 <= 0;
				CLK_64Hz <= NOT CLK_64Hz;
			 END IF;
	 END IF;
  END PROCESS;
  
  PROCESS(CLK_64Hz)
  BEGIN
    IF (CLK_64Hz'EVENT AND CLK_64Hz='0') THEN
			 COUNT_2 <= COUNT_2+1;
			 IF (COUNT_2 = 3) THEN
			   COUNT_2 <= 0;
				CLK_8Hz <= NOT CLK_8Hz;
			 END IF;
	 END IF;
  END PROCESS;
  
  PROCESS(CLK_8Hz)
  BEGIN
    IF (CLK_8Hz'EVENT AND CLK_8Hz='0') THEN
			 COUNT_3 <= COUNT_3+1;
			 IF (COUNT_3 = 3) THEN
			   COUNT_3 <= 0;
				CLK_1Hz <= NOT CLK_1Hz;
			 END IF;
	 END IF;
  END PROCESS;


END DIVIDE_SERIAL;