LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY GREENMEMEORY IS
  PORT(
  MODE_CONTROL:IN INTEGER RANGE 0 TO 7;
  COUNT_IN:IN INTEGER RANGE 0 TO 7;
  MEMORY_OUT:BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END ENTITY GREENMEMEORY;
ARCHITECTURE BEHAVE OF GREENMEMEORY IS
BEGIN
  PROCESS(couNT_IN)
  BEGIN
  END PROCESS;
END BEHAVE;