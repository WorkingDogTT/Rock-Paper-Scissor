LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--USE WORK.DIVIDER.ALL;
--USE WORK.USER1.ALL;
--USE WORK.USER2.ALL;
--USE WORK.JUDGEMENT.ALL;
--USE WORK.DISSEG.ALL;
--USE WORK.LIGHTARRAY.ALL;
--USE WORK.BTN_ARRAY.ALL;

ENTITY S1P1 IS
  PORT(
  CLK_IN:IN STD_LOGIC
  );
END ENTITY  S1P1;
ARCHITECTURE BEHAVE OF S1P1 IS
BEGIN
  PROCESS(CLK_IN)
  BEGIN
  END PROCESS;
END BEHAVE;





 
 



