LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DIVIDER IS
  PORT(
    F_1KHZ:BUFFER STD_LOGIC;
	 F_512HZ:BUFFER STD_LOGIC;
	 F_256HZ:BUFFER STD_LOGIC;
	 F_128HZ:BUFFER STD_LOGIC;
	 F_64HZ:BUFFER STD_LOGIC;
	 F_32HZ:BUFFER STD_LOGIC;
	 F_16HZ:BUFFER STD_LOGIC;
	 F_8HZ:BUFFER STD_LOGIC;
	 F_4HZ:BUFFER STD_LOGIC;
	 F_2HZ:BUFFER STD_LOGIC;
	 F_1HZ:BUFFER STD_LOGIC;
	 CLK_IN:IN STD_LOGIC
  );
END ENTITY DIVIDER;
ARCHITECTURE BEHAVE OF DIVIDER IS
BEGIN
  PROCESS(F_1KHZ)
  BEGIN
    IF CLK_IN'EVENT AND CLK_IN ='0' THEN
	    F_512HZ <= NOT F_512HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_512HZ)
  BEGIN
    IF F_512HZ'EVENT AND F_512HZ ='0' THEN
	    F_256HZ <= NOT F_256HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_256HZ)
  BEGIN
    IF F_256HZ'EVENT AND F_256HZ='0' THEN
	    F_128HZ <= NOT F_128HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_128HZ)
  BEGIN
    IF F_128HZ'EVENT AND F_128HZ='0' THEN
	    F_64HZ <= NOT F_64HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_64HZ)
  BEGIN
    IF F_64HZ'EVENT AND F_64HZ='0' THEN
	    F_32HZ <= NOT F_32HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_32HZ)
  BEGIN
    IF F_32HZ'EVENT AND F_32HZ='0' THEN
	    F_16HZ <= NOT F_16HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_16HZ)
  BEGIN
    IF F_16HZ'EVENT AND F_16HZ='0' THEN
	    F_8HZ <= NOT F_8HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_8HZ)
  BEGIN
    IF F_8HZ'EVENT AND F_8HZ='0' THEN
	    F_4HZ <= NOT F_4HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_4HZ)
  BEGIN
    IF F_4HZ'EVENT AND F_4HZ='0' THEN
	    F_2HZ <= NOT F_2HZ;
	 END IF;
  END PROCESS;
  PROCESS(F_2HZ)
  BEGIN
    IF F_2HZ'EVENT AND F_2HZ='0' THEN
	    F_1HZ <= NOT F_1HZ;
	 END IF;
  END PROCESS;
END BEHAVE;

--LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.STD_LOGIC_UNSIGNED.ALL;


--ENTITY DIVIDER_SERIAL IS
--  PORT(
--  CLK_IN    : IN STD_LOGIC;         --1kHz input clock
--  CLK_512Hz : BUFFER STD_LOGIC;     --2x diff
--  CLK_64Hz  : BUFFER STD_LOGIC;     --16x diff
--  CLK_8Hz   : BUFFER STD_LOGIC;     --128x diff
--  CLK_1Hz   : BUFFER STD_LOGIC      --1024x diff
--  );
--END DIVIDER_SERIAL;
--
--
--ARCHITECTURE DIVIDE_SERIAL OF DIVIDER_SERIAL IS
----SIGNAL COUNT:INTEGER;
----SIGNAL COUNT_MAX:INTEGER;
--  SIGNAL COUNT_1 : INTEGER RANGE 0 TO 3;
--  SIGNAL COUNT_2 : INTEGER RANGE 0 TO 3;
--  SIGNAL COUNT_3 : INTEGER RANGE 0 TO 3;
--  
--BEGIN
--
--  PROCESS(CLK_IN)
--  BEGIN
--    IF (CLK_IN'EVENT AND CLK_IN='0') THEN
--			 CLK_512Hz <= NOT CLK_512Hz;
--	 END IF;
--  END PROCESS; 
--  
--  PROCESS(CLK_512Hz)
--  BEGIN
--    IF (CLK_512Hz'EVENT AND CLK_512Hz='0') THEN
--			 
--			 IF (COUNT_1 = 3) THEN
--			   COUNT_1 <= 0;
--				CLK_64Hz <= NOT CLK_64Hz;
--			 ELSE
--			   COUNT_1 <= COUNT_1+1;
--			 END IF;
--	 END IF;
--  END PROCESS;
--  
--  PROCESS(CLK_64Hz)
--  BEGIN
--    IF (CLK_64Hz'EVENT AND CLK_64Hz='0') THEN
--			 IF (COUNT_2 = 3) THEN
--			   COUNT_2 <= 0;
--				CLK_8Hz <= NOT CLK_8Hz;
--			 ELSE
--			   COUNT_2 <= COUNT_2+1;
--			 END IF;
--	 END IF;
--  END PROCESS;
--  
--  PROCESS(CLK_8Hz)
--  BEGIN
--    IF (CLK_8Hz'EVENT AND CLK_8Hz='0') THEN
--			 
--			 IF (COUNT_3 = 3) THEN
--			   COUNT_3 <= 0;
--				CLK_1Hz <= NOT CLK_1Hz;
--			 ELSE
--				COUNT_3 <= COUNT_3+1;
--			 END IF;
--	 END IF;
--  END PROCESS;
--
--
--END DIVIDE_SERIAL;