LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--行信号读值，列信号循环写0
ENTITY BTN_DETECT IS
  PORT(
	KBROW0:IN STD_LOGIC;
	KBROW1:IN STD_LOGIC;
	KBROW2:IN STD_LOGIC;
	KBROW3:IN STD_LOGIC;
	KBROW_OUT:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END ENTITY BTN_DETECT;

ARCHITECTURE DETECTION OF BTN_DETECT IS
BEGIN
  PROCESS(KBROW0)
  BEGIN
    IF KBROW0 = '1' THEN 
	    KBROW_OUT(0) <= '1';
	 ELSE
	    KBROW_OUT(0) <= '0';
	 END IF;
  END PROCESS;
  
  PROCESS(KBROW1)
  BEGIN
    IF KBROW1 = '1' THEN 
	    KBROW_OUT(1) <= '1';
	 ELSE
	    KBROW_OUT(1) <= '0';
	 END IF;
  END PROCESS;
  
  PROCESS(KBROW2)
  BEGIN
    IF KBROW2 = '1' THEN 
	    KBROW_OUT(2) <= '1';
	 ELSE
	    KBROW_OUT(2) <= '0';
	 END IF;
  END PROCESS;
  
  PROCESS(KBROW3)
  BEGIN
    IF KBROW3 = '1' THEN 
	    KBROW_OUT(3) <= '1';
	 ELSE
	    KBROW_OUT(3) <= '0';
	 END IF;
  END PROCESS;
END DETECTION;
