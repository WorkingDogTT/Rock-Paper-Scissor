LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY USER2 IS
  PORT(
  USER2_EN:IN STD_LOGIC;
  USER2_SEL_IN:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
  USER2_SEL_OUT:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END ENTITY USER2;

ARCHITECTURE FUN OF USER2 IS
BEGIN
  PROCESS(USER2_EN,USER2_SEL_IN)
  BEGIN
    IF USER2_EN = '1' THEN
	    CASE USER2_SEL_IN IS
		   --WHEN "0000" => USER2_SLE_OUT <= "0000";  --初始化值单独出去
			WHEN "1000" => USER2_SEL_OUT <= "1000";    --石头
			WHEN "0100" => USER2_SEL_OUT <= "0100";    --剪刀
			WHEN "0010" => USER2_SEL_OUT <= "0010";    --布
			WHEN "0001" => USER2_SEL_OUT <= "0001";    --预留
		 END CASE;
	ELSE
	  USER2_SEL_OUT <= "0000" ;
	END IF;
  END PROCESS;
END FUN;