LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
                                                    --数码管译码器
ENTITY Seg_Decoder IS
   PORT(
	  Seg_select: IN STD_LOGIC_VECTOR (3 DOWNTO 0);        --显示的段码，现实的数字
	  Seg_control: OUT STD_LOGIC_VECTOR  (7 DOWNTO 0);
	  Code_input: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	  Seg_output: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
	  );
END ENTITY Seg_Decoder;

ARCHITECTURE Decode OF Seg_Decoder IS
SIGNAL Error_Flag: STD_LOGIC;
BEGIN
  Select_Seg:PROCESS(Seg_select)
  BEGIN
    CASE Seg_select IS
	   WHEN "0000"=> Seg_control<="11111110";Error_Flag<='0';
		WHEN "0001"=> Seg_control<="11111101";Error_Flag<='0';
		WHEN "0010"=> Seg_control<="11111011";Error_Flag<='0';
		WHEN "0011"=> Seg_control<="11110111";Error_Flag<='0';
		WHEN "0100"=> Seg_control<="11101111";Error_Flag<='0';
		WHEN "0101"=> Seg_control<="11011111";Error_Flag<='0';
		WHEN "0110"=> Seg_control<="10111111";Error_Flag<='0';
		WHEN "0111"=> Seg_control<="01111111";Error_Flag<='0';
		WHEN OTHERS => Seg_control<="00000000";Error_Flag<='1';
	 END CASE;	
  END PROCESS Select_Seg;
  
  Display:PROCESS(Code_input)
  BEGIN
   IF Error_Flag='0' THEN
    CASE Code_input IS
	   WHEN "0000" => Seg_output<="1111110"; --0
		WHEN "0001" => Seg_output<="0110000"; --1
		WHEN "0010" => Seg_output<="1101101"; --2
		WHEN "0011" => Seg_output<="1111001"; --3
		WHEN "0100" => Seg_output<="0110011"; --4 
		WHEN "0101" => Seg_output<="1011011"; --5
		WHEN "0110" => Seg_output<="1011111"; --6
		WHEN "0111" => Seg_output<="1110000"; --7
		WHEN"1000" => Seg_output<="1111111"; --8
		WHEN "1001" => Seg_output<="1111011"; --9
		WHEN "1111" => Seg_output<="0000000"; --灭灯指示
		WHEN "1011" => Seg_output<="0000001"; --输出 - special symbol 1
		WHEN OTHERS => Seg_output<="0000001"; --E
	 END CASE;
	ELSE 
	  Seg_output<="1001111";                --错误输出
	END IF;
  END PROCESS Display;
END  Decode;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIS IS
  PORT(
  NUM1:IN INTEGER RANGE 0 TO 5;
  NUM2:IN INTEGER RANGE 0 TO 5;
  CLK_IN:IN STD_LOGIC;
  SEG_SEL:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
  ORI_COD_OUT:OUT INTEGER
  );
END ENTITY DIS;
ARCHITECTURE DIS_UNIT OF DIS IS
SIGNAL COUNT:INTEGER RANGE 0 TO 7;
BEGIN
  TRI:PROCESS(CLK_IN)
  BEGIN
    IF CLK_IN'EVENT AND CLK_IN = '0' THEN
	    COUNT<=COUNT+1;
	 END IF;
  END PROCESS TRI;
  
  SCAN:PROCESS(COUNT,NUM1,NUM2)
  BEGIN
    CASE COUNT IS
	   WHEN 0 => SEG_SEL<= "0000";ORI_COD_OUT <= 10;   --BLANK
		WHEN 1 => SEG_SEL<= "0001";ORI_COD_OUT <= 10; --BLANK
		WHEN 2 => SEG_SEL<= "0010";ORI_COD_OUT <= NUM1;
		WHEN 3 => SEG_SEL<= "0011";ORI_COD_OUT <= 11; --special symbol 1
		WHEN 4 => SEG_SEL<= "0100";ORI_COD_OUT <= NUM2;
		WHEN 5 => SEG_SEL<= "0101";ORI_COD_OUT <= 10; --BLANK
		WHEN 6 => SEG_SEL<= "0110";ORI_COD_OUT <= 10; --BLANK
		WHEN 7 => SEG_SEL<= "0111";ORI_COD_OUT <= 10; --BLANK
		WHEN OTHERS => SEG_SEL <= "1100"; ORI_COD_OUT <= 99;--ERROR OUTPUT
	 END CASE;
  END PROCESS SCAN;  
END DIS_UNIT;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONVERTER IS
  PORT(
  ORI_COD_IN:IN INTEGER;
  COD_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END ENTITY CONVERTER;
ARCHITECTURE CONVERT OF CONVERTER IS
BEGIN
  PROCESS(ORI_COD_IN)
  BEGIN
    CASE ORI_COD_IN IS
	   WHEN 0 => COD_OUT <= "0000";
		WHEN 1 => COD_OUT <= "0001";
		WHEN 2 => COD_OUT <= "0010";
		WHEN 3 => COD_OUT <= "0011";
		WHEN 4 => COD_OUT <= "0100";
		WHEN 5 => COD_OUT <= "0101";
		WHEN 6 => COD_OUT <= "0110";
		WHEN 7 => COD_OUT <= "0111";
		WHEN 8 => COD_OUT <= "1000";
		WHEN 9 => COD_OUT <= "1001";
		WHEN 10 => COD_OUT <= "1111";
		WHEN 11 => COD_OUT <= "1011";
	   WHEN OTHERS => COD_OUT <= "1110";
	 END CASE;
  END PROCESS;
END CONVERT;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--USE WORK.DIVIDER.ALL;

ENTITY SEG_DIS IS 
  PORT(
  CLK_IN:IN STD_LOGIC;
  NUM1_IN:IN INTEGER RANGE 0 TO 5;
  NUM2_IN:IN INTEGER RANGE 0 TO 5;
  SEG_CONTROL:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  SEG_DISPLAY:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END ENTITY SEG_DIS;
ARCHITECTURE MAIN OF SEG_DIS IS 
  COMPONENT DIVIDER
     PORT(
     CLK_IN:IN STD_LOGIC;
     CLK_OUT:BUFFER STD_LOGIC;
     FRE_SET:IN INTEGER        --设置频率，必须赋给初值，单位是百Hz，否则进入默认分频状态100HZ
     );
  END COMPONENT; 
  COMPONENT CONVERTER
    PORT(
    ORI_COD_IN:IN INTEGER;
    COD_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
  END COMPONENT;
  
  COMPONENT DIS
    PORT(
    NUM1:IN INTEGER RANGE 0 TO 5;
    NUM2:IN INTEGER RANGE 0 TO 5;
    CLK_IN:IN STD_LOGIC;
    SEG_SEL:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    ORI_COD_OUT:OUT INTEGER
    );
  END COMPONENT;
  
  COMPONENT SEG_DECODER
     PORT(
	  Seg_select: IN STD_LOGIC_VECTOR (3 DOWNTO 0);       
	  Seg_control: OUT STD_LOGIC_VECTOR  (7 DOWNTO 0);
	  Code_input: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	  Seg_output: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
	  );
  END COMPONENT;
SIGNAL CLK_BUS:STD_LOGIC;
SIGNAL COD_BUFFER:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ORI_COD_BUFFER:INTEGER;
SIGNAL SEG_BUFFER:STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
  U0_divider:DIVIDER
    PORT MAP(
    CLK_IN => CLK_IN,
    CLK_OUT => CLK_BUS,
    FRE_SET => 200          --200百HZ 20KHZ
    );
  U1_converter:CONVERTER
    PORT MAP(
    ORI_COD_IN => ORI_COD_BUFFER,
    COD_OUT => COD_BUFFER
    );
  U2_DIS:DIS
    PORT MAP(
    NUM1 => NUM1_IN,
    NUM2 => NUM2_IN,
    CLK_IN => CLK_BUS,
    SEG_SEL => SEG_BUFFER,
    ORI_COD_OUT => ORI_COD_BUFFER
    );
  U3_SEG_DIS:SEG_DECODER
    PORT MAP(
	 Seg_select => SEG_BUFFER,
	 Seg_control => SEG_CONTROL,
	 Code_input => COD_BUFFER,
	 Seg_output => SEG_DISPLAY
	 );
END MAIN;
