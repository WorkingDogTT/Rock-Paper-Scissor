LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY COUNTER IS
  PORT(
  CLK_IN:IN STD_LOGIC;
  EN_IN:IN STD_LOGIC;
  STATE_OUT:BUFFER STD_LOGIC
  );
END ENTITY COUNTER;

ARCHITECTURE BEHAVE OF COUNTER IS
SIGNAL COUNT:INTEGER;
SIGNAL COUNT_MAX:INTEGER;
BEGIN
  PROCESS(CLK_IN)
  BEGIN
    IF CLK_IN'EVENT AND CLK_IN='0' THEN
	    IF EN_IN='1' THEN
		    IF COUNT>=COUNT_MAX THEN
			    STATE_OUT<='1';
			 ELSE
			    COUNT<=COUNT+1;
			 END IF;
		 ELSE
		    STATE_OUT<='0';
			 COUNT<=0;
		 END IF;
	 END IF;
  END PROCESS;
END BEHAVE;