LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REDMEMORY IS
  PORT(
  U1_MODE_CONTROL:IN INTEGER RANGE 0 TO 3;     --这里接收USER1的选择输入
  U2_MODE_CONTROL:IN INTEGER RANGE 0 TO 3;     --这里接收USER2的选择输入
  COUNT_IN:IN INTEGER RANGE 0 TO 7;            --这里接收8X8点阵的行扫数据
  MEMORY_OUT:BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0)  --输出当前的列向量
  );
END ENTITY REDMEMORY;
ARCHITECTURE BEHAVE OF REDMEMORY IS
--石头的显存定义
CONSTANT U1_R_RC_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_RC_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_RC_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="11100000";
CONSTANT U1_R_RC_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="11100000";
CONSTANT U1_R_RC_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="11100000";
CONSTANT U1_R_RC_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_RC_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_RC_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--剪刀的显存定义
CONSTANT U1_R_SC_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_SC_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_SC_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="00100000";
CONSTANT U1_R_SC_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="11000000";
CONSTANT U1_R_SC_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="11000000";
CONSTANT U1_R_SC_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="00100000";
CONSTANT U1_R_SC_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_SC_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--布的显存定义
CONSTANT U1_R_PA_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_PA_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_PA_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="01000000";
CONSTANT U1_R_PA_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="11100000";
CONSTANT U1_R_PA_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="11100000";
CONSTANT U1_R_PA_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="01000000";
CONSTANT U1_R_PA_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U1_R_PA_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--石头的显存定义
CONSTANT U2_R_RC_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_RC_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_RC_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000111";
CONSTANT U2_R_RC_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000111";
CONSTANT U2_R_RC_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000111";
CONSTANT U2_R_RC_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_RC_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_RC_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--剪刀的显存定义
CONSTANT U2_R_SC_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_SC_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_SC_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000100";
CONSTANT U2_R_SC_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000011";
CONSTANT U2_R_SC_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000011";
CONSTANT U2_R_SC_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000100";
CONSTANT U2_R_SC_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_SC_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--布的显存定义
CONSTANT U2_R_PA_R0:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_PA_R1:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_PA_R2:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000010";
CONSTANT U2_R_PA_R3:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000111";
CONSTANT U2_R_PA_R4:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000111";
CONSTANT U2_R_PA_R5:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000010";
CONSTANT U2_R_PA_R6:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
CONSTANT U2_R_PA_R7:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
--临时的显存空间
SIGNAL TEMP:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL TEMP_MOD:INTEGER RANGE 0 TO 8;
BEGIN
  PROCESS(U1_MODE_CONTROL,U2_MODE_CONTROL)
  BEGIN
     CASE U1_MODE_CONTROL IS
	    WHEN 0 => 
		   CASE U2_MODE_CONTROL IS
			    WHEN 0 => 
				   TEMP_MOD <= 0;   --Rock against Rock
				 WHEN 1 =>
				   TEMP_MOD <= 1;   --Rock against Scissor
             WHEN 2 =>
				   TEMP_MOD <= 2;   --Rock against Paper
				 WHEN OTHERS => 	
			END CASE;
		 WHEN 1 => 
		 	 CASE U2_MODE_CONTROL IS
			    WHEN 0 => 
				   TEMP_MOD <= 3;   --Scissor against Rock
				 WHEN 1 =>
				   TEMP_MOD <= 4;   --Scissor against Scissor
             WHEN 2 =>
				   TEMP_MOD <= 5;   --Scissor against Paper
				 WHEN OTHERS => 	
			END CASE;
		 WHEN 2 => 
		 	  CASE U2_MODE_CONTROL IS
			    WHEN 0 => 
				   TEMP_MOD <= 6;   --Paper against Rock
				 WHEN 1 =>
				   TEMP_MOD <= 7;   --Paper against Scissor
             WHEN 2 =>
				   TEMP_MOD <= 8;   --Paper against Paper 
		       WHEN OTHERS => 
		     END CASE;
	    WHEN OTHERS => 
	  END CASE;
  END PROCESS;
  
  PROCESS(COUNT_IN,TEMP_MOD)
  BEGIN
    CASE COUNT_IN IS
	   WHEN 0 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R0 OR U2_R_RC_R0;
			 WHEN 1 => TEMP <= U1_R_RC_R0 OR U2_R_SC_R0;
			 WHEN 2 => TEMP <= U1_R_RC_R0 OR U2_R_PA_R0;
			 WHEN 3 => TEMP <= U1_R_SC_R0 OR U2_R_RC_R0;
			 WHEN 4 => TEMP <= U1_R_SC_R0 OR U2_R_SC_R0;
			 WHEN 5 => TEMP <= U1_R_SC_R0 OR U2_R_PA_R0;
			 WHEN 6 => TEMP <= U1_R_PA_R0 OR U2_R_RC_R0;
			 WHEN 7 => TEMP <= U1_R_PA_R0 OR U2_R_SC_R0;
			 WHEN 8 => TEMP <= U1_R_PA_R0 OR U2_R_PA_R0;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 1 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R1 OR U2_R_RC_R1;
			 WHEN 1 => TEMP <= U1_R_RC_R1 OR U2_R_SC_R1;
			 WHEN 2 => TEMP <= U1_R_RC_R1 OR U2_R_PA_R1;
			 WHEN 3 => TEMP <= U1_R_SC_R1 OR U2_R_RC_R1;
			 WHEN 4 => TEMP <= U1_R_SC_R1 OR U2_R_SC_R1;
			 WHEN 5 => TEMP <= U1_R_SC_R1 OR U2_R_PA_R1;
			 WHEN 6 => TEMP <= U1_R_PA_R1 OR U2_R_RC_R1;
			 WHEN 7 => TEMP <= U1_R_PA_R1 OR U2_R_SC_R1;
			 WHEN 8 => TEMP <= U1_R_PA_R1 OR U2_R_PA_R1;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 2 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R2 OR U2_R_RC_R2;
			 WHEN 1 => TEMP <= U1_R_RC_R2 OR U2_R_SC_R2;
			 WHEN 2 => TEMP <= U1_R_RC_R2 OR U2_R_PA_R2;
			 WHEN 3 => TEMP <= U1_R_SC_R2 OR U2_R_RC_R2;
			 WHEN 4 => TEMP <= U1_R_SC_R2 OR U2_R_SC_R2;
			 WHEN 5 => TEMP <= U1_R_SC_R2 OR U2_R_PA_R2;
			 WHEN 6 => TEMP <= U1_R_PA_R2 OR U2_R_RC_R2;
			 WHEN 7 => TEMP <= U1_R_PA_R2 OR U2_R_SC_R2;
			 WHEN 8 => TEMP <= U1_R_PA_R2 OR U2_R_PA_R2;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 3 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R3 OR U2_R_RC_R3;
			 WHEN 1 => TEMP <= U1_R_RC_R3 OR U2_R_SC_R3;
			 WHEN 2 => TEMP <= U1_R_RC_R3 OR U2_R_PA_R3;
			 WHEN 3 => TEMP <= U1_R_SC_R3 OR U2_R_RC_R3;
			 WHEN 4 => TEMP <= U1_R_SC_R3 OR U2_R_SC_R3;
			 WHEN 5 => TEMP <= U1_R_SC_R3 OR U2_R_PA_R3;
			 WHEN 6 => TEMP <= U1_R_PA_R3 OR U2_R_RC_R3;
			 WHEN 7 => TEMP <= U1_R_PA_R3 OR U2_R_SC_R3;
			 WHEN 8 => TEMP <= U1_R_PA_R3 OR U2_R_PA_R3;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 4 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R4 OR U2_R_RC_R4;
			 WHEN 1 => TEMP <= U1_R_RC_R4 OR U2_R_SC_R4;
			 WHEN 2 => TEMP <= U1_R_RC_R4 OR U2_R_PA_R4;
			 WHEN 3 => TEMP <= U1_R_SC_R4 OR U2_R_RC_R4;
			 WHEN 4 => TEMP <= U1_R_SC_R4 OR U2_R_SC_R4;
			 WHEN 5 => TEMP <= U1_R_SC_R4 OR U2_R_PA_R4;
			 WHEN 6 => TEMP <= U1_R_PA_R4 OR U2_R_RC_R4;
			 WHEN 7 => TEMP <= U1_R_PA_R4 OR U2_R_SC_R4;
			 WHEN 8 => TEMP <= U1_R_PA_R4 OR U2_R_PA_R4;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 5 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R5 OR U2_R_RC_R5;
			 WHEN 1 => TEMP <= U1_R_RC_R5 OR U2_R_SC_R5;
			 WHEN 2 => TEMP <= U1_R_RC_R5 OR U2_R_PA_R5;
			 WHEN 3 => TEMP <= U1_R_SC_R5 OR U2_R_RC_R5;
			 WHEN 4 => TEMP <= U1_R_SC_R5 OR U2_R_SC_R5;
			 WHEN 5 => TEMP <= U1_R_SC_R5 OR U2_R_PA_R5;
			 WHEN 6 => TEMP <= U1_R_PA_R5 OR U2_R_RC_R5;
			 WHEN 7 => TEMP <= U1_R_PA_R5 OR U2_R_SC_R5;
			 WHEN 8 => TEMP <= U1_R_PA_R5 OR U2_R_PA_R5;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 6 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R6 OR U2_R_RC_R6;
			 WHEN 1 => TEMP <= U1_R_RC_R6 OR U2_R_SC_R6;
			 WHEN 2 => TEMP <= U1_R_RC_R6 OR U2_R_PA_R6;
			 WHEN 3 => TEMP <= U1_R_SC_R6 OR U2_R_RC_R6;
			 WHEN 4 => TEMP <= U1_R_SC_R6 OR U2_R_SC_R6;
			 WHEN 5 => TEMP <= U1_R_SC_R6 OR U2_R_PA_R6;
			 WHEN 6 => TEMP <= U1_R_PA_R6 OR U2_R_RC_R6;
			 WHEN 7 => TEMP <= U1_R_PA_R6 OR U2_R_SC_R6;
			 WHEN 8 => TEMP <= U1_R_PA_R6 OR U2_R_PA_R6;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN 7 =>
		  CASE TEMP_MOD IS
		    WHEN 0 => TEMP <= U1_R_RC_R7 OR U2_R_RC_R7;
			 WHEN 1 => TEMP <= U1_R_RC_R7 OR U2_R_SC_R7;
			 WHEN 2 => TEMP <= U1_R_RC_R7 OR U2_R_PA_R7;
			 WHEN 3 => TEMP <= U1_R_SC_R7 OR U2_R_RC_R7;
			 WHEN 4 => TEMP <= U1_R_SC_R7 OR U2_R_SC_R7;
			 WHEN 5 => TEMP <= U1_R_SC_R7 OR U2_R_PA_R7;
			 WHEN 6 => TEMP <= U1_R_PA_R7 OR U2_R_RC_R7;
			 WHEN 7 => TEMP <= U1_R_PA_R7 OR U2_R_SC_R7;
			 WHEN 8 => TEMP <= U1_R_PA_R7 OR U2_R_PA_R7;
			 WHEN OTHERS =>  TEMP <= "00000000";
		  END CASE;
		WHEN OTHERS =>
	 END CASE;
  END PROCESS;
  
  PROCESS(TEMP)
  BEGIN
    MEMORY_OUT <= TEMP;
  END PROCESS;
END BEHAVE; 